`timescale 1ns / 1ps
module datapath(input  logic        clk, reset,
                input  logic        memtoreg, pcsrc,
                input  logic        alusrc, regdst,
                input  logic        regwrite, jump,
                input  logic [2:0]  alucontrol,
                output logic        zero,
                output logic [31:0] pc,
                input  logic [31:0] instr,
                output logic [31:0] aluout, writedata,
                input  logic [31:0] readdata,
                input  logic        shift,    // added
                output logic        sign,     // added
                input  logic        li,       // added
                input  logic        zfr       // added
                );

  logic [4:0]  writereg;
  logic [31:0] pcnext, pcnextbr, pcplus4, pcbranch;
  logic [31:0] signimm, signimmsh;
  logic [31:0] RD1, RD2;        // added for clarity
  logic [31:0] srca, srcb;
  logic [31:0] liout;       // added
  logic [31:0] result;
  logic [31:0] zfrout;      // added
  
  // debug displayer
  always_comb begin
      //$display("shift: %b", shift);
      //$display("li: %b, liout: %h, aluout: %h", li, liout, aluout);
      $display("dataaddr: %h, writedata: %h", aluout, RD2);
  end

  // next PC logic
  flopr #(32) pcreg(clk, reset, pcnext, pc);
  adder #(32) pcadd1(pc, 32'b100, 'b0, pcplus4); //So we adjust this to use the more complex adder; wmt-modification
  sl2         immsh(signimm, signimmsh);
  adder #(32) pcadd2(pcplus4, signimmsh, 'b0, pcbranch); //See comment above
  mux2 #(32)  pcbrmux(pcplus4, pcbranch, pcsrc, pcnextbr);
  mux2 #(32)  pcmux(pcnextbr, {pcplus4[31:28], 
                    instr[25:0], 2'b00}, jump, pcnext);

  // register file logic
  assign    writedata = RD2;    //added
  regfile     rf(clk, regwrite, instr[25:21], instr[20:16], 
                 writereg, result, RD1, RD2); // modded srca to RD1, writedata to RD2
  mux2 #(5)   wrmux(instr[20:16], instr[15:11],
                    regdst, writereg);
  mux2 #(32)  limux(aluout, {16'b0, instr[15:0]}, li, liout);   // added for li
  mux2 #(32)  resmux(liout, readdata, memtoreg, result);        // aluout to liout
  signext     se(instr[15:0], signimm);

  // ALU logic
  // addded srcamux for sll, zero-extend 5-bit shamt to 32-bits
  // added zfrmux for zfr, bit mask generated by 0xFFFF_FFFE << RD2[4:0]
  mux2 #(32)  srcamux(RD1, {27'b0, instr[10:6]}, shift, srca);
  mux2 #(32)  srcbmux(RD2, signimm, alusrc, srcb);
  mux2 #(32)  zfrmux(srcb, 32'hFFFF_FFFE << RD2[4:0], zfr, zfrout); // added for zfr
  alu         alu(srca, zfrout, alucontrol, aluout, zero, sign);
  
endmodule